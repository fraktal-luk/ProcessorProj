----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:03:19 05/05/2016 
-- Design Name: 
-- Module Name:    SubunitDispatch - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

use work.ProcBasicDefs.all;
use work.Helpers.all;

use work.ProcInstructionsNew.all;

use work.NewPipelineData.all;

use work.GeneralPipeDev.all;

--use work.CommonRouting.all;
use work.TEMP_DEV.all;

use work.ProcLogicIQ.all;

use work.ProcComponents.all;


entity SubunitDispatch is
	port(
		clk: in std_logic;
		reset: in std_logic;
		en: in std_logic;
		
	 	prevSending: in std_logic;
	 	nextAccepting: in std_logic;
		

	 	stageDataIn: in InstructionState;		
		acceptingOut: out std_logic;
		sendingOut: out std_logic;
		stageDataOut: out InstructionState;
		
		execEventSignal: in std_logic;
		execCausing: in InstructionState;
		intSignal: in std_logic;
		
		ai: in ArgStatusInfo;
		resultVals: in MwordArray(0 to N_RES_TAGS-1);
		regValues: in MwordArray(0 to 2);
		
		dispatchDataOut: out InstructionState
	);
end SubunitDispatch;


architecture Behavioral of SubunitDispatch is
	signal dispatchData, dispatchDataNext, dispatchDataUpdated,
				inputDataWithArgs: InstructionState := defaultInstructionState;
	signal flowDriveDispatch: FlowDriveSimple := (others=>'0');											
	signal flowResponseDispatch: FlowResponseSimple := (others=>'0');		
begin	
	acceptingOut <= flowResponseDispatch.accepting;
	flowDriveDispatch.prevSending <= prevSending;
										
	DISPATCH_SYNCHRONOUS: process(clk)
	begin
		if rising_edge(clk) then
			if en = '1' then
				dispatchData <= dispatchDataNext;
			end if;				
		end if;
	end process;
	
	inputDataWithArgs <= getDispatchArgValues(stageDataIn, resultVals);
	dispatchDataNext <= stageSimpleNext(dispatchData, --Updated, 
														inputDataWithArgs,
													flowResponseDispatch.living,
													flowResponseDispatch.sending, 
													--flowDriveDispatch.prevSending);
														flowResponseDispatch.accepting);
	dispatchDataUpdated <= updateDispatchArgs(dispatchData, resultVals, regValues, ai); 
		
	-- Don't allow exec if args somehow are not actualy ready!		
	flowDriveDispatch.lockSend <= --not asDispatch.readyAll;
							BLOCK_ISSUE_WHEN_MISSING and isNonzero(dispatchDataUpdated.argValues.missing);
	
	-- Dispatch pipe logic
	SIMPLE_SLOT_LOGIC_DISPATCH_A: SimplePipeLogic port map(
		clk => clk, reset => reset, en => en,
		flowDrive => flowDriveDispatch,
		flowResponse => flowResponseDispatch
	);	
		
	DISPATCH_A_KILL: block
		signal before: std_logic;
		signal a, b: std_logic_vector(7 downto 0);
	begin
		a <= execCausing.groupTag;
		b <= dispatchData.groupTag;	

		IQ_KILLER: entity work.CompareBefore8 port map(
			inA =>  a,
			inB =>  b,
			outC => before
		);
		
		--before <= '0'; --
					--tagBefore(a, b);			
		flowDriveDispatch.kill <= killByTag(before, execEventSignal, intSignal);
										-- before and execEventSignal; 	
	end block;			
				
	stageDataOut <= dispatchDataUpdated;
	sendingOut <= flowResponseDispatch.sending;

	flowDriveDispatch.nextAccepting <= nextAccepting;
	
	dispatchDataOut <= dispatchData;
end Behavioral;


architecture Alternative of SubunitDispatch is
	signal stageDataM, stageDataStored: StageDataMulti := DEFAULT_STAGE_DATA_MULTI;
	signal inputDataWithArgs, dispatchDataUpdated:
					InstructionState := defaultInstructionState;
		signal lockSend: std_logic := '0';
begin

	inputDataWithArgs <= getDispatchArgValues(stageDataIn, resultVals);

	stageDataM.fullMask(0) <= prevSending;
	stageDataM.data(0) <= inputDataWithArgs;
	
	BASIC_LOGIC: entity work.GenericStageMulti(SingleTagged)
	port map(
		clk => clk, reset => reset, en => en,
		
		prevSending => prevSending,
		nextAccepting => nextAccepting,
		
		stageDataIn => stageDataM,
		acceptingOut => acceptingOut,
		sendingOut => sendingOut,
		stageDataOut => stageDataStored,
		
		execEventSignal => execEventSignal,
		execCausing => execCausing,
		lockCommand => '0'
	);

	dispatchDataUpdated <= updateDispatchArgs(stageDataStored.data(0), resultVals, regValues, ai); 

		-- CAREFUL: this does nothing. To make it work:
		--											nextAcceptingEffective <= nextAccepting and not lockSend
		lockSend <= BLOCK_ISSUE_WHEN_MISSING and isNonzero(dispatchDataUpdated.argValues.missing);
	
	stageDataOut <= dispatchDataUpdated;
	
end Alternative;


